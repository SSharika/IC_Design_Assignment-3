module adder (
    input a,
    input b,
    output reg sum
);

always@*


 sum = a + b;

endmodule

